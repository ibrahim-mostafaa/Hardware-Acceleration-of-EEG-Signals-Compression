module xor_1bit (
input wire a,b,
output wire y); 

assign y = a^b; 
endmodule 